`timescale 1ns/1ps
module pes_elevator_tb;

reg [7:0]request_floor;
reg [7:0]in_current_floor;
reg clk;
reg reset;
reg over_time;
reg over_weight;

wire direction;
wire complete;
wire door_alert;
wire weight_alert;
wire [7:0] out_current_floor;

pes_elevator UUT(
.request_floor (request_floor),
.in_current_floor (in_current_floor),
.clk(clk),
.reset (reset),
.direction (direction),
.out_current_floor (out_current_floor),
.complete (complete),
.over_time (over_time),
.over_weight (over_weight),
.door_alert (door_alert),
.weight_alert (weight_alert));



//Generate the clock and test the circuit with different inputs
initial
begin
  $dumpfile ("pes_elevator_tb.vcd"); 
  $dumpvars(0,pes_elevatorr_tb);
#0 clk =1'b0; reset =1'b0; over_time=1'b0; over_weight=1'b0;
//#50 reset =1'b0;
#25 request_floor = 8'b00000001; in_current_floor = 8'b10000000;
#25 reset =1;
#50 reset =0;

#50 over_time =1;
#50 over_time =0;
//#50 reset =1'b1;
//#70 reset =1'b0;
#50 over_weight =1;
#100 over_weight =0;

//#50 reset = 1'b1;
#300 $finish;
end
always
#25 clk=~clk;

endmodule


